<svg width="161" height="219" viewBox="0 0 161 219" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M46.7441 1.29456C46.7441 1.29456 23.6367 14.8036 14.3434 29.3158C0.941181 50.2443 -0.270035 68.4576 3.07349 93.865C8.12843 132.277 19.0869 154.206 58.5214 171.924C97.9558 189.643 120.065 199.576 159.5 217.295" stroke="white" stroke-width="3"/>
</svg>
